
module debug_subsystem (
	clk_clk,
	cpu_debug_bus_bridge_0_interrupt_irq,
	ppu_debug_bus_bridge_0_interrupt_irq,
	reset_reset_n,
	to_external_bus_bridge_0_external_interface_acknowledge,
	to_external_bus_bridge_0_external_interface_irq,
	to_external_bus_bridge_0_external_interface_address,
	to_external_bus_bridge_0_external_interface_bus_enable,
	to_external_bus_bridge_0_external_interface_byte_enable,
	to_external_bus_bridge_0_external_interface_rw,
	to_external_bus_bridge_0_external_interface_write_data,
	to_external_bus_bridge_0_external_interface_read_data,
	to_external_bus_bridge_1_external_interface_acknowledge,
	to_external_bus_bridge_1_external_interface_irq,
	to_external_bus_bridge_1_external_interface_address,
	to_external_bus_bridge_1_external_interface_bus_enable,
	to_external_bus_bridge_1_external_interface_byte_enable,
	to_external_bus_bridge_1_external_interface_rw,
	to_external_bus_bridge_1_external_interface_write_data,
	to_external_bus_bridge_1_external_interface_read_data,
	clk_1_clk_clk,
	clk_1_clk_reset_reset_n,
	clk_ppu_0_clk_clk,
	clk_ppu_0_clk_reset_reset_n);	

	input		clk_clk;
	output		cpu_debug_bus_bridge_0_interrupt_irq;
	output		ppu_debug_bus_bridge_0_interrupt_irq;
	input		reset_reset_n;
	input		to_external_bus_bridge_0_external_interface_acknowledge;
	input		to_external_bus_bridge_0_external_interface_irq;
	output	[15:0]	to_external_bus_bridge_0_external_interface_address;
	output		to_external_bus_bridge_0_external_interface_bus_enable;
	output	[1:0]	to_external_bus_bridge_0_external_interface_byte_enable;
	output		to_external_bus_bridge_0_external_interface_rw;
	output	[15:0]	to_external_bus_bridge_0_external_interface_write_data;
	input	[15:0]	to_external_bus_bridge_0_external_interface_read_data;
	input		to_external_bus_bridge_1_external_interface_acknowledge;
	input		to_external_bus_bridge_1_external_interface_irq;
	output	[15:0]	to_external_bus_bridge_1_external_interface_address;
	output		to_external_bus_bridge_1_external_interface_bus_enable;
	output	[1:0]	to_external_bus_bridge_1_external_interface_byte_enable;
	output		to_external_bus_bridge_1_external_interface_rw;
	output	[15:0]	to_external_bus_bridge_1_external_interface_write_data;
	input	[15:0]	to_external_bus_bridge_1_external_interface_read_data;
	output		clk_1_clk_clk;
	output		clk_1_clk_reset_reset_n;
	output		clk_ppu_0_clk_clk;
	output		clk_ppu_0_clk_reset_reset_n;
endmodule
