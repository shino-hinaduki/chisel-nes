// debug_subsystem.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module debug_subsystem (
		input  wire        clk_clk,                                                 //                                         clk.clk
		output wire        clk_1_clk_clk,                                           //                                   clk_1_clk.clk
		output wire        clk_1_clk_reset_reset_n,                                 //                             clk_1_clk_reset.reset_n
		output wire        clk_ppu_0_clk_clk,                                       //                               clk_ppu_0_clk.clk
		output wire        clk_ppu_0_clk_reset_reset_n,                             //                         clk_ppu_0_clk_reset.reset_n
		output wire        cpu_debug_bus_bridge_0_interrupt_irq,                    //            cpu_debug_bus_bridge_0_interrupt.irq
		output wire        ppu_debug_bus_bridge_0_interrupt_irq,                    //            ppu_debug_bus_bridge_0_interrupt.irq
		input  wire        reset_reset_n,                                           //                                       reset.reset_n
		input  wire        to_external_bus_bridge_0_external_interface_acknowledge, // to_external_bus_bridge_0_external_interface.acknowledge
		input  wire        to_external_bus_bridge_0_external_interface_irq,         //                                            .irq
		output wire [15:0] to_external_bus_bridge_0_external_interface_address,     //                                            .address
		output wire        to_external_bus_bridge_0_external_interface_bus_enable,  //                                            .bus_enable
		output wire [1:0]  to_external_bus_bridge_0_external_interface_byte_enable, //                                            .byte_enable
		output wire        to_external_bus_bridge_0_external_interface_rw,          //                                            .rw
		output wire [15:0] to_external_bus_bridge_0_external_interface_write_data,  //                                            .write_data
		input  wire [15:0] to_external_bus_bridge_0_external_interface_read_data,   //                                            .read_data
		input  wire        to_external_bus_bridge_1_external_interface_acknowledge, // to_external_bus_bridge_1_external_interface.acknowledge
		input  wire        to_external_bus_bridge_1_external_interface_irq,         //                                            .irq
		output wire [15:0] to_external_bus_bridge_1_external_interface_address,     //                                            .address
		output wire        to_external_bus_bridge_1_external_interface_bus_enable,  //                                            .bus_enable
		output wire [1:0]  to_external_bus_bridge_1_external_interface_byte_enable, //                                            .byte_enable
		output wire        to_external_bus_bridge_1_external_interface_rw,          //                                            .rw
		output wire [15:0] to_external_bus_bridge_1_external_interface_write_data,  //                                            .write_data
		input  wire [15:0] to_external_bus_bridge_1_external_interface_read_data    //                                            .read_data
	);

	wire         pll_0_outclk1_clk;                                                 // pll_0:outclk_1 -> [mm_interconnect_1:pll_0_outclk1_clk, mm_interconnect_2:pll_0_outclk1_clk, ppu_clock_bridge_0:s0_clk, ppu_debug_bus_bridge_0:clk, rst_controller_003:clk, rst_controller_004:clk]
	wire         cpu_clock_bridge_0_m0_waitrequest;                                 // mm_interconnect_0:cpu_clock_bridge_0_m0_waitrequest -> cpu_clock_bridge_0:m0_waitrequest
	wire  [31:0] cpu_clock_bridge_0_m0_readdata;                                    // mm_interconnect_0:cpu_clock_bridge_0_m0_readdata -> cpu_clock_bridge_0:m0_readdata
	wire         cpu_clock_bridge_0_m0_debugaccess;                                 // cpu_clock_bridge_0:m0_debugaccess -> mm_interconnect_0:cpu_clock_bridge_0_m0_debugaccess
	wire  [15:0] cpu_clock_bridge_0_m0_address;                                     // cpu_clock_bridge_0:m0_address -> mm_interconnect_0:cpu_clock_bridge_0_m0_address
	wire         cpu_clock_bridge_0_m0_read;                                        // cpu_clock_bridge_0:m0_read -> mm_interconnect_0:cpu_clock_bridge_0_m0_read
	wire   [3:0] cpu_clock_bridge_0_m0_byteenable;                                  // cpu_clock_bridge_0:m0_byteenable -> mm_interconnect_0:cpu_clock_bridge_0_m0_byteenable
	wire         cpu_clock_bridge_0_m0_readdatavalid;                               // mm_interconnect_0:cpu_clock_bridge_0_m0_readdatavalid -> cpu_clock_bridge_0:m0_readdatavalid
	wire  [31:0] cpu_clock_bridge_0_m0_writedata;                                   // cpu_clock_bridge_0:m0_writedata -> mm_interconnect_0:cpu_clock_bridge_0_m0_writedata
	wire         cpu_clock_bridge_0_m0_write;                                       // cpu_clock_bridge_0:m0_write -> mm_interconnect_0:cpu_clock_bridge_0_m0_write
	wire   [0:0] cpu_clock_bridge_0_m0_burstcount;                                  // cpu_clock_bridge_0:m0_burstcount -> mm_interconnect_0:cpu_clock_bridge_0_m0_burstcount
	wire         mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_chipselect;  // mm_interconnect_0:cpu_debug_bus_bridge_0_avalon_slave_chipselect -> cpu_debug_bus_bridge_0:avalon_chipselect
	wire  [15:0] mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_readdata;    // cpu_debug_bus_bridge_0:avalon_readdata -> mm_interconnect_0:cpu_debug_bus_bridge_0_avalon_slave_readdata
	wire         mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_waitrequest; // cpu_debug_bus_bridge_0:avalon_waitrequest -> mm_interconnect_0:cpu_debug_bus_bridge_0_avalon_slave_waitrequest
	wire  [14:0] mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_address;     // mm_interconnect_0:cpu_debug_bus_bridge_0_avalon_slave_address -> cpu_debug_bus_bridge_0:avalon_address
	wire         mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_read;        // mm_interconnect_0:cpu_debug_bus_bridge_0_avalon_slave_read -> cpu_debug_bus_bridge_0:avalon_read
	wire   [1:0] mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_byteenable;  // mm_interconnect_0:cpu_debug_bus_bridge_0_avalon_slave_byteenable -> cpu_debug_bus_bridge_0:avalon_byteenable
	wire         mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_write;       // mm_interconnect_0:cpu_debug_bus_bridge_0_avalon_slave_write -> cpu_debug_bus_bridge_0:avalon_write
	wire  [15:0] mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_writedata;   // mm_interconnect_0:cpu_debug_bus_bridge_0_avalon_slave_writedata -> cpu_debug_bus_bridge_0:avalon_writedata
	wire         ppu_clock_bridge_0_m0_waitrequest;                                 // mm_interconnect_1:ppu_clock_bridge_0_m0_waitrequest -> ppu_clock_bridge_0:m0_waitrequest
	wire  [31:0] ppu_clock_bridge_0_m0_readdata;                                    // mm_interconnect_1:ppu_clock_bridge_0_m0_readdata -> ppu_clock_bridge_0:m0_readdata
	wire         ppu_clock_bridge_0_m0_debugaccess;                                 // ppu_clock_bridge_0:m0_debugaccess -> mm_interconnect_1:ppu_clock_bridge_0_m0_debugaccess
	wire  [15:0] ppu_clock_bridge_0_m0_address;                                     // ppu_clock_bridge_0:m0_address -> mm_interconnect_1:ppu_clock_bridge_0_m0_address
	wire         ppu_clock_bridge_0_m0_read;                                        // ppu_clock_bridge_0:m0_read -> mm_interconnect_1:ppu_clock_bridge_0_m0_read
	wire   [3:0] ppu_clock_bridge_0_m0_byteenable;                                  // ppu_clock_bridge_0:m0_byteenable -> mm_interconnect_1:ppu_clock_bridge_0_m0_byteenable
	wire         ppu_clock_bridge_0_m0_readdatavalid;                               // mm_interconnect_1:ppu_clock_bridge_0_m0_readdatavalid -> ppu_clock_bridge_0:m0_readdatavalid
	wire  [31:0] ppu_clock_bridge_0_m0_writedata;                                   // ppu_clock_bridge_0:m0_writedata -> mm_interconnect_1:ppu_clock_bridge_0_m0_writedata
	wire         ppu_clock_bridge_0_m0_write;                                       // ppu_clock_bridge_0:m0_write -> mm_interconnect_1:ppu_clock_bridge_0_m0_write
	wire   [0:0] ppu_clock_bridge_0_m0_burstcount;                                  // ppu_clock_bridge_0:m0_burstcount -> mm_interconnect_1:ppu_clock_bridge_0_m0_burstcount
	wire         mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_chipselect;  // mm_interconnect_1:ppu_debug_bus_bridge_0_avalon_slave_chipselect -> ppu_debug_bus_bridge_0:avalon_chipselect
	wire  [15:0] mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_readdata;    // ppu_debug_bus_bridge_0:avalon_readdata -> mm_interconnect_1:ppu_debug_bus_bridge_0_avalon_slave_readdata
	wire         mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_waitrequest; // ppu_debug_bus_bridge_0:avalon_waitrequest -> mm_interconnect_1:ppu_debug_bus_bridge_0_avalon_slave_waitrequest
	wire  [14:0] mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_address;     // mm_interconnect_1:ppu_debug_bus_bridge_0_avalon_slave_address -> ppu_debug_bus_bridge_0:avalon_address
	wire         mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_read;        // mm_interconnect_1:ppu_debug_bus_bridge_0_avalon_slave_read -> ppu_debug_bus_bridge_0:avalon_read
	wire   [1:0] mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_byteenable;  // mm_interconnect_1:ppu_debug_bus_bridge_0_avalon_slave_byteenable -> ppu_debug_bus_bridge_0:avalon_byteenable
	wire         mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_write;       // mm_interconnect_1:ppu_debug_bus_bridge_0_avalon_slave_write -> ppu_debug_bus_bridge_0:avalon_write
	wire  [15:0] mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_writedata;   // mm_interconnect_1:ppu_debug_bus_bridge_0_avalon_slave_writedata -> ppu_debug_bus_bridge_0:avalon_writedata
	wire  [31:0] jtag_to_avalon_master_0_master_readdata;                           // mm_interconnect_2:jtag_to_avalon_master_0_master_readdata -> jtag_to_avalon_master_0:master_readdata
	wire         jtag_to_avalon_master_0_master_waitrequest;                        // mm_interconnect_2:jtag_to_avalon_master_0_master_waitrequest -> jtag_to_avalon_master_0:master_waitrequest
	wire  [31:0] jtag_to_avalon_master_0_master_address;                            // jtag_to_avalon_master_0:master_address -> mm_interconnect_2:jtag_to_avalon_master_0_master_address
	wire         jtag_to_avalon_master_0_master_read;                               // jtag_to_avalon_master_0:master_read -> mm_interconnect_2:jtag_to_avalon_master_0_master_read
	wire   [3:0] jtag_to_avalon_master_0_master_byteenable;                         // jtag_to_avalon_master_0:master_byteenable -> mm_interconnect_2:jtag_to_avalon_master_0_master_byteenable
	wire         jtag_to_avalon_master_0_master_readdatavalid;                      // mm_interconnect_2:jtag_to_avalon_master_0_master_readdatavalid -> jtag_to_avalon_master_0:master_readdatavalid
	wire         jtag_to_avalon_master_0_master_write;                              // jtag_to_avalon_master_0:master_write -> mm_interconnect_2:jtag_to_avalon_master_0_master_write
	wire  [31:0] jtag_to_avalon_master_0_master_writedata;                          // jtag_to_avalon_master_0:master_writedata -> mm_interconnect_2:jtag_to_avalon_master_0_master_writedata
	wire  [31:0] mm_interconnect_2_sysid_0_control_slave_readdata;                  // sysid_0:readdata -> mm_interconnect_2:sysid_0_control_slave_readdata
	wire   [0:0] mm_interconnect_2_sysid_0_control_slave_address;                   // mm_interconnect_2:sysid_0_control_slave_address -> sysid_0:address
	wire  [31:0] mm_interconnect_2_cpu_clock_bridge_0_s0_readdata;                  // cpu_clock_bridge_0:s0_readdata -> mm_interconnect_2:cpu_clock_bridge_0_s0_readdata
	wire         mm_interconnect_2_cpu_clock_bridge_0_s0_waitrequest;               // cpu_clock_bridge_0:s0_waitrequest -> mm_interconnect_2:cpu_clock_bridge_0_s0_waitrequest
	wire         mm_interconnect_2_cpu_clock_bridge_0_s0_debugaccess;               // mm_interconnect_2:cpu_clock_bridge_0_s0_debugaccess -> cpu_clock_bridge_0:s0_debugaccess
	wire  [15:0] mm_interconnect_2_cpu_clock_bridge_0_s0_address;                   // mm_interconnect_2:cpu_clock_bridge_0_s0_address -> cpu_clock_bridge_0:s0_address
	wire         mm_interconnect_2_cpu_clock_bridge_0_s0_read;                      // mm_interconnect_2:cpu_clock_bridge_0_s0_read -> cpu_clock_bridge_0:s0_read
	wire   [3:0] mm_interconnect_2_cpu_clock_bridge_0_s0_byteenable;                // mm_interconnect_2:cpu_clock_bridge_0_s0_byteenable -> cpu_clock_bridge_0:s0_byteenable
	wire         mm_interconnect_2_cpu_clock_bridge_0_s0_readdatavalid;             // cpu_clock_bridge_0:s0_readdatavalid -> mm_interconnect_2:cpu_clock_bridge_0_s0_readdatavalid
	wire         mm_interconnect_2_cpu_clock_bridge_0_s0_write;                     // mm_interconnect_2:cpu_clock_bridge_0_s0_write -> cpu_clock_bridge_0:s0_write
	wire  [31:0] mm_interconnect_2_cpu_clock_bridge_0_s0_writedata;                 // mm_interconnect_2:cpu_clock_bridge_0_s0_writedata -> cpu_clock_bridge_0:s0_writedata
	wire   [0:0] mm_interconnect_2_cpu_clock_bridge_0_s0_burstcount;                // mm_interconnect_2:cpu_clock_bridge_0_s0_burstcount -> cpu_clock_bridge_0:s0_burstcount
	wire  [31:0] mm_interconnect_2_ppu_clock_bridge_0_s0_readdata;                  // ppu_clock_bridge_0:s0_readdata -> mm_interconnect_2:ppu_clock_bridge_0_s0_readdata
	wire         mm_interconnect_2_ppu_clock_bridge_0_s0_waitrequest;               // ppu_clock_bridge_0:s0_waitrequest -> mm_interconnect_2:ppu_clock_bridge_0_s0_waitrequest
	wire         mm_interconnect_2_ppu_clock_bridge_0_s0_debugaccess;               // mm_interconnect_2:ppu_clock_bridge_0_s0_debugaccess -> ppu_clock_bridge_0:s0_debugaccess
	wire  [15:0] mm_interconnect_2_ppu_clock_bridge_0_s0_address;                   // mm_interconnect_2:ppu_clock_bridge_0_s0_address -> ppu_clock_bridge_0:s0_address
	wire         mm_interconnect_2_ppu_clock_bridge_0_s0_read;                      // mm_interconnect_2:ppu_clock_bridge_0_s0_read -> ppu_clock_bridge_0:s0_read
	wire   [3:0] mm_interconnect_2_ppu_clock_bridge_0_s0_byteenable;                // mm_interconnect_2:ppu_clock_bridge_0_s0_byteenable -> ppu_clock_bridge_0:s0_byteenable
	wire         mm_interconnect_2_ppu_clock_bridge_0_s0_readdatavalid;             // ppu_clock_bridge_0:s0_readdatavalid -> mm_interconnect_2:ppu_clock_bridge_0_s0_readdatavalid
	wire         mm_interconnect_2_ppu_clock_bridge_0_s0_write;                     // mm_interconnect_2:ppu_clock_bridge_0_s0_write -> ppu_clock_bridge_0:s0_write
	wire  [31:0] mm_interconnect_2_ppu_clock_bridge_0_s0_writedata;                 // mm_interconnect_2:ppu_clock_bridge_0_s0_writedata -> ppu_clock_bridge_0:s0_writedata
	wire   [0:0] mm_interconnect_2_ppu_clock_bridge_0_s0_burstcount;                // mm_interconnect_2:ppu_clock_bridge_0_s0_burstcount -> ppu_clock_bridge_0:s0_burstcount
	wire         rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [cpu_clock_bridge_0:m0_reset, mm_interconnect_0:cpu_clock_bridge_0_m0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ppu_clock_bridge_0_m0_reset_reset_bridge_in_reset_reset, ppu_clock_bridge_0:m0_reset]
	wire         jtag_to_avalon_master_0_master_reset_reset;                        // jtag_to_avalon_master_0:master_reset_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_003:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                // rst_controller_001:reset_out -> [cpu_clock_bridge_0:s0_reset, mm_interconnect_2:cpu_clock_bridge_0_s0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                                // rst_controller_002:reset_out -> [cpu_debug_bus_bridge_0:reset, mm_interconnect_0:cpu_debug_bus_bridge_0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_003_reset_out_reset;                                // rst_controller_003:reset_out -> [mm_interconnect_2:ppu_clock_bridge_0_s0_reset_reset_bridge_in_reset_reset, ppu_clock_bridge_0:s0_reset]
	wire         rst_controller_004_reset_out_reset;                                // rst_controller_004:reset_out -> [mm_interconnect_1:ppu_debug_bus_bridge_0_reset_reset_bridge_in_reset_reset, ppu_debug_bus_bridge_0:reset]
	wire         rst_controller_005_reset_out_reset;                                // rst_controller_005:reset_out -> [mm_interconnect_2:jtag_to_avalon_master_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:sysid_0_reset_reset_bridge_in_reset_reset, sysid_0:reset_n]

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (16),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) cpu_clock_bridge_0 (
		.m0_clk           (clk_clk),                                               //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),                        // m0_reset.reset
		.s0_clk           (clk_1_clk_clk),                                         //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                    // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_2_cpu_clock_bridge_0_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_2_cpu_clock_bridge_0_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_2_cpu_clock_bridge_0_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_2_cpu_clock_bridge_0_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_2_cpu_clock_bridge_0_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_2_cpu_clock_bridge_0_s0_address),       //         .address
		.s0_write         (mm_interconnect_2_cpu_clock_bridge_0_s0_write),         //         .write
		.s0_read          (mm_interconnect_2_cpu_clock_bridge_0_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_2_cpu_clock_bridge_0_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_2_cpu_clock_bridge_0_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (cpu_clock_bridge_0_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (cpu_clock_bridge_0_m0_readdata),                        //         .readdata
		.m0_readdatavalid (cpu_clock_bridge_0_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (cpu_clock_bridge_0_m0_burstcount),                      //         .burstcount
		.m0_writedata     (cpu_clock_bridge_0_m0_writedata),                       //         .writedata
		.m0_address       (cpu_clock_bridge_0_m0_address),                         //         .address
		.m0_write         (cpu_clock_bridge_0_m0_write),                           //         .write
		.m0_read          (cpu_clock_bridge_0_m0_read),                            //         .read
		.m0_byteenable    (cpu_clock_bridge_0_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (cpu_clock_bridge_0_m0_debugaccess)                      //         .debugaccess
	);

	debug_subsystem_cpu_debug_bus_bridge_0 cpu_debug_bus_bridge_0 (
		.clk                (clk_1_clk_clk),                                                     //                clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                //              reset.reset
		.avalon_address     (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_address),     //       avalon_slave.address
		.avalon_byteenable  (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_byteenable),  //                   .byteenable
		.avalon_chipselect  (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_chipselect),  //                   .chipselect
		.avalon_read        (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_read),        //                   .read
		.avalon_write       (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_write),       //                   .write
		.avalon_writedata   (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_writedata),   //                   .writedata
		.avalon_readdata    (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_readdata),    //                   .readdata
		.avalon_waitrequest (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_waitrequest), //                   .waitrequest
		.avalon_irq         (cpu_debug_bus_bridge_0_interrupt_irq),                              //          interrupt.irq
		.acknowledge        (to_external_bus_bridge_0_external_interface_acknowledge),           // external_interface.export
		.irq                (to_external_bus_bridge_0_external_interface_irq),                   //                   .export
		.address            (to_external_bus_bridge_0_external_interface_address),               //                   .export
		.bus_enable         (to_external_bus_bridge_0_external_interface_bus_enable),            //                   .export
		.byte_enable        (to_external_bus_bridge_0_external_interface_byte_enable),           //                   .export
		.rw                 (to_external_bus_bridge_0_external_interface_rw),                    //                   .export
		.write_data         (to_external_bus_bridge_0_external_interface_write_data),            //                   .export
		.read_data          (to_external_bus_bridge_0_external_interface_read_data)              //                   .export
	);

	debug_subsystem_jtag_to_avalon_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_to_avalon_master_0 (
		.clk_clk              (clk_clk),                                      //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                               //    clk_reset.reset
		.master_address       (jtag_to_avalon_master_0_master_address),       //       master.address
		.master_readdata      (jtag_to_avalon_master_0_master_readdata),      //             .readdata
		.master_read          (jtag_to_avalon_master_0_master_read),          //             .read
		.master_write         (jtag_to_avalon_master_0_master_write),         //             .write
		.master_writedata     (jtag_to_avalon_master_0_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_to_avalon_master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_to_avalon_master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_to_avalon_master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   (jtag_to_avalon_master_0_master_reset_reset)    // master_reset.reset
	);

	debug_subsystem_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (clk_1_clk_clk),     // outclk0.clk
		.outclk_1 (pll_0_outclk1_clk), // outclk1.clk
		.locked   ()                   // (terminated)
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (16),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) ppu_clock_bridge_0 (
		.m0_clk           (clk_clk),                                               //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),                        // m0_reset.reset
		.s0_clk           (pll_0_outclk1_clk),                                     //   s0_clk.clk
		.s0_reset         (rst_controller_003_reset_out_reset),                    // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_2_ppu_clock_bridge_0_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_2_ppu_clock_bridge_0_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_2_ppu_clock_bridge_0_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_2_ppu_clock_bridge_0_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_2_ppu_clock_bridge_0_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_2_ppu_clock_bridge_0_s0_address),       //         .address
		.s0_write         (mm_interconnect_2_ppu_clock_bridge_0_s0_write),         //         .write
		.s0_read          (mm_interconnect_2_ppu_clock_bridge_0_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_2_ppu_clock_bridge_0_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_2_ppu_clock_bridge_0_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (ppu_clock_bridge_0_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (ppu_clock_bridge_0_m0_readdata),                        //         .readdata
		.m0_readdatavalid (ppu_clock_bridge_0_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (ppu_clock_bridge_0_m0_burstcount),                      //         .burstcount
		.m0_writedata     (ppu_clock_bridge_0_m0_writedata),                       //         .writedata
		.m0_address       (ppu_clock_bridge_0_m0_address),                         //         .address
		.m0_write         (ppu_clock_bridge_0_m0_write),                           //         .write
		.m0_read          (ppu_clock_bridge_0_m0_read),                            //         .read
		.m0_byteenable    (ppu_clock_bridge_0_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (ppu_clock_bridge_0_m0_debugaccess)                      //         .debugaccess
	);

	debug_subsystem_ppu_debug_bus_bridge_0 ppu_debug_bus_bridge_0 (
		.clk                (pll_0_outclk1_clk),                                                 //                clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                //              reset.reset
		.avalon_address     (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_address),     //       avalon_slave.address
		.avalon_byteenable  (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_byteenable),  //                   .byteenable
		.avalon_chipselect  (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_chipselect),  //                   .chipselect
		.avalon_read        (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_read),        //                   .read
		.avalon_write       (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_write),       //                   .write
		.avalon_writedata   (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_writedata),   //                   .writedata
		.avalon_readdata    (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_readdata),    //                   .readdata
		.avalon_waitrequest (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_waitrequest), //                   .waitrequest
		.avalon_irq         (ppu_debug_bus_bridge_0_interrupt_irq),                              //          interrupt.irq
		.acknowledge        (to_external_bus_bridge_1_external_interface_acknowledge),           // external_interface.export
		.irq                (to_external_bus_bridge_1_external_interface_irq),                   //                   .export
		.address            (to_external_bus_bridge_1_external_interface_address),               //                   .export
		.bus_enable         (to_external_bus_bridge_1_external_interface_bus_enable),            //                   .export
		.byte_enable        (to_external_bus_bridge_1_external_interface_byte_enable),           //                   .export
		.rw                 (to_external_bus_bridge_1_external_interface_rw),                    //                   .export
		.write_data         (to_external_bus_bridge_1_external_interface_write_data),            //                   .export
		.read_data          (to_external_bus_bridge_1_external_interface_read_data)              //                   .export
	);

	debug_subsystem_sysid_0 sysid_0 (
		.clock    (clk_clk),                                          //           clk.clk
		.reset_n  (~rst_controller_005_reset_out_reset),              //         reset.reset_n
		.readdata (mm_interconnect_2_sysid_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_2_sysid_0_control_slave_address)   //              .address
	);

	debug_subsystem_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                            (clk_clk),                                                           //                                          clk_0_clk.clk
		.pll_0_outclk0_clk                                        (clk_1_clk_clk),                                                     //                                      pll_0_outclk0.clk
		.cpu_clock_bridge_0_m0_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                                    //  cpu_clock_bridge_0_m0_reset_reset_bridge_in_reset.reset
		.cpu_debug_bus_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                // cpu_debug_bus_bridge_0_reset_reset_bridge_in_reset.reset
		.cpu_clock_bridge_0_m0_address                            (cpu_clock_bridge_0_m0_address),                                     //                              cpu_clock_bridge_0_m0.address
		.cpu_clock_bridge_0_m0_waitrequest                        (cpu_clock_bridge_0_m0_waitrequest),                                 //                                                   .waitrequest
		.cpu_clock_bridge_0_m0_burstcount                         (cpu_clock_bridge_0_m0_burstcount),                                  //                                                   .burstcount
		.cpu_clock_bridge_0_m0_byteenable                         (cpu_clock_bridge_0_m0_byteenable),                                  //                                                   .byteenable
		.cpu_clock_bridge_0_m0_read                               (cpu_clock_bridge_0_m0_read),                                        //                                                   .read
		.cpu_clock_bridge_0_m0_readdata                           (cpu_clock_bridge_0_m0_readdata),                                    //                                                   .readdata
		.cpu_clock_bridge_0_m0_readdatavalid                      (cpu_clock_bridge_0_m0_readdatavalid),                               //                                                   .readdatavalid
		.cpu_clock_bridge_0_m0_write                              (cpu_clock_bridge_0_m0_write),                                       //                                                   .write
		.cpu_clock_bridge_0_m0_writedata                          (cpu_clock_bridge_0_m0_writedata),                                   //                                                   .writedata
		.cpu_clock_bridge_0_m0_debugaccess                        (cpu_clock_bridge_0_m0_debugaccess),                                 //                                                   .debugaccess
		.cpu_debug_bus_bridge_0_avalon_slave_address              (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_address),     //                cpu_debug_bus_bridge_0_avalon_slave.address
		.cpu_debug_bus_bridge_0_avalon_slave_write                (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_write),       //                                                   .write
		.cpu_debug_bus_bridge_0_avalon_slave_read                 (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_read),        //                                                   .read
		.cpu_debug_bus_bridge_0_avalon_slave_readdata             (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_readdata),    //                                                   .readdata
		.cpu_debug_bus_bridge_0_avalon_slave_writedata            (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_writedata),   //                                                   .writedata
		.cpu_debug_bus_bridge_0_avalon_slave_byteenable           (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_byteenable),  //                                                   .byteenable
		.cpu_debug_bus_bridge_0_avalon_slave_waitrequest          (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_waitrequest), //                                                   .waitrequest
		.cpu_debug_bus_bridge_0_avalon_slave_chipselect           (mm_interconnect_0_cpu_debug_bus_bridge_0_avalon_slave_chipselect)   //                                                   .chipselect
	);

	debug_subsystem_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                            (clk_clk),                                                           //                                          clk_0_clk.clk
		.pll_0_outclk1_clk                                        (pll_0_outclk1_clk),                                                 //                                      pll_0_outclk1.clk
		.ppu_clock_bridge_0_m0_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                                    //  ppu_clock_bridge_0_m0_reset_reset_bridge_in_reset.reset
		.ppu_debug_bus_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                                // ppu_debug_bus_bridge_0_reset_reset_bridge_in_reset.reset
		.ppu_clock_bridge_0_m0_address                            (ppu_clock_bridge_0_m0_address),                                     //                              ppu_clock_bridge_0_m0.address
		.ppu_clock_bridge_0_m0_waitrequest                        (ppu_clock_bridge_0_m0_waitrequest),                                 //                                                   .waitrequest
		.ppu_clock_bridge_0_m0_burstcount                         (ppu_clock_bridge_0_m0_burstcount),                                  //                                                   .burstcount
		.ppu_clock_bridge_0_m0_byteenable                         (ppu_clock_bridge_0_m0_byteenable),                                  //                                                   .byteenable
		.ppu_clock_bridge_0_m0_read                               (ppu_clock_bridge_0_m0_read),                                        //                                                   .read
		.ppu_clock_bridge_0_m0_readdata                           (ppu_clock_bridge_0_m0_readdata),                                    //                                                   .readdata
		.ppu_clock_bridge_0_m0_readdatavalid                      (ppu_clock_bridge_0_m0_readdatavalid),                               //                                                   .readdatavalid
		.ppu_clock_bridge_0_m0_write                              (ppu_clock_bridge_0_m0_write),                                       //                                                   .write
		.ppu_clock_bridge_0_m0_writedata                          (ppu_clock_bridge_0_m0_writedata),                                   //                                                   .writedata
		.ppu_clock_bridge_0_m0_debugaccess                        (ppu_clock_bridge_0_m0_debugaccess),                                 //                                                   .debugaccess
		.ppu_debug_bus_bridge_0_avalon_slave_address              (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_address),     //                ppu_debug_bus_bridge_0_avalon_slave.address
		.ppu_debug_bus_bridge_0_avalon_slave_write                (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_write),       //                                                   .write
		.ppu_debug_bus_bridge_0_avalon_slave_read                 (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_read),        //                                                   .read
		.ppu_debug_bus_bridge_0_avalon_slave_readdata             (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_readdata),    //                                                   .readdata
		.ppu_debug_bus_bridge_0_avalon_slave_writedata            (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_writedata),   //                                                   .writedata
		.ppu_debug_bus_bridge_0_avalon_slave_byteenable           (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_byteenable),  //                                                   .byteenable
		.ppu_debug_bus_bridge_0_avalon_slave_waitrequest          (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_waitrequest), //                                                   .waitrequest
		.ppu_debug_bus_bridge_0_avalon_slave_chipselect           (mm_interconnect_1_ppu_debug_bus_bridge_0_avalon_slave_chipselect)   //                                                   .chipselect
	);

	debug_subsystem_mm_interconnect_2 mm_interconnect_2 (
		.clk_0_clk_clk                                                 (clk_clk),                                               //                                               clk_0_clk.clk
		.pll_0_outclk0_clk                                             (clk_1_clk_clk),                                         //                                           pll_0_outclk0.clk
		.pll_0_outclk1_clk                                             (pll_0_outclk1_clk),                                     //                                           pll_0_outclk1.clk
		.cpu_clock_bridge_0_s0_reset_reset_bridge_in_reset_reset       (rst_controller_001_reset_out_reset),                    //       cpu_clock_bridge_0_s0_reset_reset_bridge_in_reset.reset
		.jtag_to_avalon_master_0_clk_reset_reset_bridge_in_reset_reset (rst_controller_005_reset_out_reset),                    // jtag_to_avalon_master_0_clk_reset_reset_bridge_in_reset.reset
		.ppu_clock_bridge_0_s0_reset_reset_bridge_in_reset_reset       (rst_controller_003_reset_out_reset),                    //       ppu_clock_bridge_0_s0_reset_reset_bridge_in_reset.reset
		.sysid_0_reset_reset_bridge_in_reset_reset                     (rst_controller_005_reset_out_reset),                    //                     sysid_0_reset_reset_bridge_in_reset.reset
		.jtag_to_avalon_master_0_master_address                        (jtag_to_avalon_master_0_master_address),                //                          jtag_to_avalon_master_0_master.address
		.jtag_to_avalon_master_0_master_waitrequest                    (jtag_to_avalon_master_0_master_waitrequest),            //                                                        .waitrequest
		.jtag_to_avalon_master_0_master_byteenable                     (jtag_to_avalon_master_0_master_byteenable),             //                                                        .byteenable
		.jtag_to_avalon_master_0_master_read                           (jtag_to_avalon_master_0_master_read),                   //                                                        .read
		.jtag_to_avalon_master_0_master_readdata                       (jtag_to_avalon_master_0_master_readdata),               //                                                        .readdata
		.jtag_to_avalon_master_0_master_readdatavalid                  (jtag_to_avalon_master_0_master_readdatavalid),          //                                                        .readdatavalid
		.jtag_to_avalon_master_0_master_write                          (jtag_to_avalon_master_0_master_write),                  //                                                        .write
		.jtag_to_avalon_master_0_master_writedata                      (jtag_to_avalon_master_0_master_writedata),              //                                                        .writedata
		.cpu_clock_bridge_0_s0_address                                 (mm_interconnect_2_cpu_clock_bridge_0_s0_address),       //                                   cpu_clock_bridge_0_s0.address
		.cpu_clock_bridge_0_s0_write                                   (mm_interconnect_2_cpu_clock_bridge_0_s0_write),         //                                                        .write
		.cpu_clock_bridge_0_s0_read                                    (mm_interconnect_2_cpu_clock_bridge_0_s0_read),          //                                                        .read
		.cpu_clock_bridge_0_s0_readdata                                (mm_interconnect_2_cpu_clock_bridge_0_s0_readdata),      //                                                        .readdata
		.cpu_clock_bridge_0_s0_writedata                               (mm_interconnect_2_cpu_clock_bridge_0_s0_writedata),     //                                                        .writedata
		.cpu_clock_bridge_0_s0_burstcount                              (mm_interconnect_2_cpu_clock_bridge_0_s0_burstcount),    //                                                        .burstcount
		.cpu_clock_bridge_0_s0_byteenable                              (mm_interconnect_2_cpu_clock_bridge_0_s0_byteenable),    //                                                        .byteenable
		.cpu_clock_bridge_0_s0_readdatavalid                           (mm_interconnect_2_cpu_clock_bridge_0_s0_readdatavalid), //                                                        .readdatavalid
		.cpu_clock_bridge_0_s0_waitrequest                             (mm_interconnect_2_cpu_clock_bridge_0_s0_waitrequest),   //                                                        .waitrequest
		.cpu_clock_bridge_0_s0_debugaccess                             (mm_interconnect_2_cpu_clock_bridge_0_s0_debugaccess),   //                                                        .debugaccess
		.ppu_clock_bridge_0_s0_address                                 (mm_interconnect_2_ppu_clock_bridge_0_s0_address),       //                                   ppu_clock_bridge_0_s0.address
		.ppu_clock_bridge_0_s0_write                                   (mm_interconnect_2_ppu_clock_bridge_0_s0_write),         //                                                        .write
		.ppu_clock_bridge_0_s0_read                                    (mm_interconnect_2_ppu_clock_bridge_0_s0_read),          //                                                        .read
		.ppu_clock_bridge_0_s0_readdata                                (mm_interconnect_2_ppu_clock_bridge_0_s0_readdata),      //                                                        .readdata
		.ppu_clock_bridge_0_s0_writedata                               (mm_interconnect_2_ppu_clock_bridge_0_s0_writedata),     //                                                        .writedata
		.ppu_clock_bridge_0_s0_burstcount                              (mm_interconnect_2_ppu_clock_bridge_0_s0_burstcount),    //                                                        .burstcount
		.ppu_clock_bridge_0_s0_byteenable                              (mm_interconnect_2_ppu_clock_bridge_0_s0_byteenable),    //                                                        .byteenable
		.ppu_clock_bridge_0_s0_readdatavalid                           (mm_interconnect_2_ppu_clock_bridge_0_s0_readdatavalid), //                                                        .readdatavalid
		.ppu_clock_bridge_0_s0_waitrequest                             (mm_interconnect_2_ppu_clock_bridge_0_s0_waitrequest),   //                                                        .waitrequest
		.ppu_clock_bridge_0_s0_debugaccess                             (mm_interconnect_2_ppu_clock_bridge_0_s0_debugaccess),   //                                                        .debugaccess
		.sysid_0_control_slave_address                                 (mm_interconnect_2_sysid_0_control_slave_address),       //                                   sysid_0_control_slave.address
		.sysid_0_control_slave_readdata                                (mm_interconnect_2_sysid_0_control_slave_readdata)       //                                                        .readdata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (jtag_to_avalon_master_0_master_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (jtag_to_avalon_master_0_master_reset_reset), // reset_in1.reset
		.clk            (clk_1_clk_clk),                              //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_1_clk_clk),                      //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (jtag_to_avalon_master_0_master_reset_reset), // reset_in1.reset
		.clk            (pll_0_outclk1_clk),                          //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_0_outclk1_clk),                  //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	assign clk_ppu_0_clk_clk = clk_clk;

	assign clk_1_clk_reset_reset_n = reset_reset_n;

	assign clk_ppu_0_clk_reset_reset_n = reset_reset_n;

endmodule
